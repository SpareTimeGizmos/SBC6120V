//++
//sbc6120_ume2.v - SBC6120/V test bench for Spare Time Gizmos UME2 board
//Copyright (C) 2011-2014 by Spare Time Gizmos.  All rights reserved.
//
// DESCRIPTION:
//   This module runs the SBC6120V on the Spare Time Gizmos UME2 board, and
// the actual FPGA on this board is the Spartan 3E XC3S500-5PQ208.
//
// REVISION HISTORY:
// 27-Jan-11 RLA  new file.
//  1-Jan-14  RLA  Remove global reset net.  Add initial blocks instead.
//--
//000000011111111112222222222333333333344444444445555555555666666666677777777778
//345678901234567890123456789012345678901234567890123456789012345678901234567890
`include "sbc6120_h.v"

//   These includes are required because we have ifdefs around the instances of
// these modules.  If we don't explicitly include them, Xilinx can't seem to
// figure out the module hierarchy.  XST will complain that these modules aren't
// defined, even though they're obviously part of the project ...
`include "fp6120.v"
`include "ds1302.v"
`include "cfcard.v"
`include "sdcard.v"


module ume2_clkgen
  //++
  //   This module uses one of the nifty Xilinx digital clock managers to
  // generate both a CPU clock and a VGA pixel clock.  The system clock is
  // nominally 50Mhz, and a 25MHz CPU clock is generated by using the DLL part
  // of the DCM to divide by two.  At the same time we use the frequency
  // synthesizer part of the same DCM to generate a 28MHz VGA dot clock by
  // multiplying the ratio 17/30.  That's all there is to it!
  //
  //   IMPORTANT - notice that we don't use the locked output of the DCM.  The
  // FPGA startup MUST BE CONFIGURED TO WAIT FOR DCM LOCKED!
  //--
( 
  input  clock_50mhz, 	// 50Mhz system clock
  output cpuclk, 	// 25Mhz cpu clock
  output vgaclk 	// 28Mhz VGA dot clock
);
  parameter CPU_CLOCK_DIVIDE     =  4;
  parameter PIXEL_CLOCK_MULTIPLY = 17;
  parameter PIXEL_CLOCK_DIVIDE   = 30;

  // Locals ...
  wire clkdv_unbuf;	// unbuffered DCM CLKDV (cpuclk)
  wire clkfx_unbuf;	// unbuffered DCM CLKFX (vgaclk)
  wire clk0_unbuf;	// unbuffered DCM CLK0 output
  wire clkfb_buf;	// buffered CLK0 for DCM feedback

  // Here's the magic part!
  DCM_SP #(
    .CLKDV_DIVIDE(CPU_CLOCK_DIVIDE),
    .CLKFX_DIVIDE(PIXEL_CLOCK_DIVIDE), .CLKFX_MULTIPLY(PIXEL_CLOCK_MULTIPLY),
    .CLK_FEEDBACK("1X"), .FACTORY_JF(16'h8080),
    .STARTUP_WAIT("TRUE")
   ) clkdcm (
    .CLKIN(clock_50mhz), .CLK0(clk0_unbuf), .CLKFB(clkfb_buf), 
    .CLKDV(clkdv_unbuf), .CLKFX(clkfx_unbuf), .LOCKED(),
    .DSSEN(1'b0), .PSCLK(1'b0), .PSEN(1'b0), .PSINCDEC(1'b0), .RST(1'b0)
  );
  
  //   Buffer all the clocks we generate with global buffers, and that includes
  // sticking a BUFG in the feedback path for the DCM.  That's so the DCM will
  // automatically compensate for the 1ns or so delay added by the BUFG.  This
  // application is not very critical and that's overkill, but it's the "right" 
  // way to do it...
  BUFG cpuclk_bufg    (.I(clkdv_unbuf), .O(cpuclk));
  BUFG vgaclk_bufg    (.I(clkfx_unbuf), .O(vgaclk));
  BUFG clkdcm_fb_bufg (.I(clk0_unbuf),  .O(clkfb_buf));
endmodule // ume2_clkgen


module ume2_beeper (
  //++
  //   This module drives the piezo beeper on the UME2, and when triggered
  // it generates a fixed length tone of about 6kHz for 300ms.  Note that this
  // is driven by the VGA clock - it's connected to the VT52, so it's convenient
  // to have it exist in that clock domain - and the timing is based on the
  // 28.322MHz VGA dot clock.
  //--
  input  clock,			// free running 50Mhz system clock
  input  enable, 		// asserted for one tick to trigger the bell
  output speaker, 		// push-pull speaker drive output
  output speaker_n		//  ...
);
  parameter LOG2_DELAY = 23; 	// about 300ms delay at 28.322MHz
  parameter MAX_DELAY = 2**LOG2_DELAY-1;
  reg [LOG2_DELAY-1:0] count;	// bell timer
  initial count = 0;		// the initial state is "bell off"!

  // When triggered, just count down from MAX_DELAY to zero ...  
  always @(posedge clock)
    if (enable)
      count <= 2**LOG2_DELAY-1;
    else if (count != 0)
      count <= count-1;

  //   The two speaker outputs toggle, out of phase, as long as the count is
  // non-zero.  We cheat and just use one of the bits int he counter to toggle
  // the outputs - this gives a frequency of about 6kHz and saves us from
  // needing yet another counter.
  assign speaker   = (count != 0) ?  count[13] : 0;
  assign speaker_n = (count != 0) ? ~count[13] : 0;
endmodule // ume2_beeper


module ume2_scanner
  //++
  //   This module generates the column drive for the UME2 seven segment
  // displays and keypad.  These three devices (two six digit LED displays and
  // a 4x4 keypad) share the same column drive and so their interfaces have to
  // be coordinated.  The column drive is just a simple barrel shifter that
  // rotates a single zero bit, the column drives being active low, thru the
  // six scan outputs.  We also produce a key_tick output that signals the 
  // keypad logic that it's time to sample the key state. 
  //--
#(
  parameter CLOCK_FREQUENCY = 50_000_000,
  parameter SCAN_FREQUENCY =       1_500
) (
  input 	   clock,	// free running 50Mhz system clock
  output reg [5:0] scan_n,	// 7 segment LEDs and keypad column drive
  output           key_tick	// tells the keypad when to sample the keys
);
  // Generate a 1.5kHz scan clock ...
  wire scan_tick;
  ck_divider #(.IN_FREQ(CLOCK_FREQUENCY), .OUT_FREQ(SCAN_FREQUENCY))
    scan_clock (.clock(clock), .out(scan_tick));

  //   A subtle point is that key_tick is an asynchronous output, so it will
  // actually become true in the same clock cycle where scan_tick is asserted.
  // The scan_n outputs, however, are registered so they won't actually change
  // until the next clock cycle _after_ the one where scan_tick was asserted.
  // That means key_tick will preceed the columns changing by one clock, which
  // is exactly what we want to happen.
  assign key_tick = scan_tick;

  // The scan register always as 5 ones and exactly one zero ...
  initial scan_n = 6'b111110;
  
  // Now we can generate the column drive ....
  always @(posedge clock)
    if (scan_tick) scan_n <= {scan_n[4:0], scan_n[5]};
endmodule // ume2_scanner


module ume2_display
  //++
  //   This module drives the UME2 seven segment LED displays.  There are two
  // such displays with six digits each, and the data for them is specified as
  // two 24 bit vectors with four bits of BCD data per digit.  The column drive
  // for the displays is generated separately by the ume2_scanner module, and
  // this module is purely combinatorial.  It's basically just a seven segment
  // decoder and multiplexor.
  //
  //   If the ALLOW_HEX parameter is defined as 1, then the four BCD bits for
  // each digit are decoded with a hex font (or as close as you can come to
  // such a thing on a seven segment display).  If ALLOW_HEX is zero then the
  // digits are decoded with a decimal font and the BCD values A..F generate
  // special characters -
  //
  //	A - TBA (blanked for now)
  //	B - TBA (blanked for now)
  //	C - TBA (blanked for now)
  //	D - TBA (blanked for now)
  //	E - "-"
  //	F - blank
  //--
#(
  parameter ALLOW_HEX = 0
) (
  output [6:0] 	adisp,		// address (upper) 7 segment LEDs segment drive
  output [6:0] 	ddisp,		// data    (lower) "   "   "   "   "   "    "
  input  [5:0] 	scan_n,		// column drive from ume2_scanner module
  input  [23:0]	addr,		// data for the address displays
  input  [23:0]	data		//  "    "   "  data     "   "
);

  // This function decodes BCD to seven segments ...
  function [6:0] decode (input [3:0] bcd);
  begin
    case (bcd)
      4'h0: decode =             7'b0111111;		   // 0
      4'h1: decode =             7'b0000110;		   // 1
      4'h2: decode =             7'b1011011;		   // 2
      4'h3: decode =             7'b1001111;		   // 3
      4'h4: decode =             7'b1100110;		   // 4
      4'h5: decode =             7'b1101101;		   // 5
      4'h6: decode =             7'b1111101;		   // 6
      4'h7: decode =             7'b0000111;		   // 7
      4'h8: decode =             7'b1111111;		   // 8
      4'h9: decode =             7'b1101111;		   // 9
      4'hA: decode = ALLOW_HEX ? 7'b1110111 : 7'b0000000;  // A
      4'hB: decode = ALLOW_HEX ? 7'b1111100 : 7'b0000000;  // b
      4'hC: decode = ALLOW_HEX ? 7'b0111001 : 7'b0000000;  // C
      4'hD: decode = ALLOW_HEX ? 7'b1011110 : 7'b0000000;  // d
      4'hE: decode = ALLOW_HEX ? 7'b1111001 : 7'b1000000;  // E
      4'hF: decode = ALLOW_HEX ? 7'b1110001 : 7'b0000000;  // F
    endcase // case (bcd)
  end
  endfunction // decode

  // Two muxes to select the correct BCD digit from the input vectors ...
  reg [3:0] a_bcd, d_bcd;
  always @* begin
    case (scan_n)
      6'b011111:  a_bcd = addr[23:20];
      6'b101111:  a_bcd = addr[19:16];
      6'b110111:  a_bcd = addr[15:12];
      6'b111011:  a_bcd = addr[11: 8];
      6'b111101:  a_bcd = addr[ 7: 4];
      6'b111110:  a_bcd = addr[ 3: 0];
      default:    a_bcd = 0; 
    endcase // case (scan_n)
  end
  always @* begin
    case (scan_n)
      6'b011111:  d_bcd = data[23:20];
      6'b101111:  d_bcd = data[19:16];
      6'b110111:  d_bcd = data[15:12];
      6'b111011:  d_bcd = data[11: 8];
      6'b111101:  d_bcd = data[ 7: 4];
      6'b111110:  d_bcd = data[ 3: 0];
      default:    d_bcd = 0; 
    endcase // case (scan_n)
  end

  // And two seven segment decoders to drive the display ...
  assign adisp = decode(a_bcd);
  assign ddisp = decode(d_bcd);
endmodule // ume2_display


// UME2 keypad definitions for the SBC6120...
//   BTW, the actual mapping of the 16 bit raw key code to the positions on
// the keypad goes like this -
//
//               col 1     col 2    col 3     col 4
//             --------  --------  --------  --------
//    row 1  | 16'h1000  16'h2000  16'h4000  16'h8000
//    row 2  | 16'h0100  16'h0200  16'h0400  16'h0800
//    row 3  | 16'h0010  16'h0020  16'h0040  16'h0080
//    row 4  | 16'h0001  16'h0002  16'h0004  16'h0008
`define KEY_0		16'h0001
`define KEY_1		16'h0002
`define KEY_2		16'h0010
`define KEY_3		16'h0020
`define KEY_4		16'h0100
`define KEY_5		16'h0200
`define KEY_6		16'h1000
`define KEY_7		16'h2000
`define KEY_LA		16'h4000
`define KEY_LXA		16'h8000
`define KEY_EXAM	16'h0400
`define KEY_DEP		16'h0800
`define KEY_CLEAR	16'h0040
`define KEY_CONT	16'h0080
`define KEY_BOOT	16'h0008
// The rest are shifted keys ...
`define KEY_SHIFT	16'h0004
`define KEY_POST	(`KEY_SHIFT | `KEY_7)
`define KEY_MQ		(`KEY_SHIFT | `KEY_3)
`define KEY_AC		(`KEY_SHIFT | `KEY_2)
`define KEY_FLAGS	(`KEY_SHIFT | `KEY_1)
`define KEY_MD		(`KEY_SHIFT | `KEY_0)


module ume2_keypad
  //++
  //   This module scans the 4x4 matrix UME2 keypad and outputs a simple 16
  // bit vector corresponding to the key(s) pressed.  A key_press strobe is
  // asserted for one clock tick every time a new key is pressed, but there
  // is no strobe or other indication when a key is released.  The keyboard
  // is debounced by keeping a running record of the last four samples, and
  // no action is taken until all four samples agree.  With a scan clock of
  // 1.5kHz, that gives a debounce time of about 16ms.
  //
  //   Note that the keypad rows are our inputs, and the keypad columns are
  // shared with the seven segment LED columns.  That means that we don't get
  // to drive the column outputs - they're generated by the ume2_scanner
  // module and shared by both this module and ume2_display.  
  //--
(
  input             clock,	// free running 50Mhz system clock
  input      [5:0]  scan_n,	// keypad column drive
  input             key_tick,	// timing tick to sample keypad state
  input      [3:0]  keyrow_n,	// keypad row inputs
  output reg [15:0] keys,	// hex value of key currently pressed
  output reg        key_press	// one tick "key pressed" strobe
);
  // Locals ...
  reg [15:0] rawkeys, key0, key1, key2, key3;

  // The keyrow inputs are asynchronous and must be synchronized first ...
  wire [3:0] keyrow_sync_n;
  synchronize_level sl0 (clock, keyrow_n[0], keyrow_sync_n[0]);
  synchronize_level sl1 (clock, keyrow_n[1], keyrow_sync_n[1]);
  synchronize_level sl2 (clock, keyrow_n[2], keyrow_sync_n[2]);
  synchronize_level sl3 (clock, keyrow_n[3], keyrow_sync_n[3]);

  // Define the initial state ...
  initial begin
    key0 = 0;  key1 = 0;  key2 = 0;  key3 = 0;
    rawkeys = 0;  keys = 0;  key_press = 0;
  end
  
  //   The keypad only has four columns (where as the LED displays have six) so
  // for the first four scan clocks we accumulate a bitmap of the keys that are
  // currently pressed.
  always @(posedge clock)
    if (key_tick & ~&scan_n[3:0])
      rawkeys <= {~keyrow_sync_n, rawkeys[15:4]};

  //   And then on the fifth scan clock we encode the keymap to a single hex
  // value and save that.  We keep the last four encoded values for debouncing
  // and pretty much ignore them until all four agree...
  always @(posedge clock)
    if (key_tick & ~scan_n[4]) begin
      key3 <= key2;  key2 <= key1;  key1 <= key0;  key0 <= rawkeys;
    end
  wire key_valid = (rawkeys==key0) & (key0==key1) & (key1==key2) & (key2==key3);

  //  The key output always holds the last valid key state detected ...
  always @(posedge clock)
    if (key_valid) keys <= key3;

  //   The problem now is to generate a key_press output that's asserted when
  // ever a new key is pressed.  It should not be asserted when a previously
  // pressed key continues to be pressed, not should it be asserted when a
  // key is released.  The latter is true even if there are also other keys
  // pressed at the same time.  Sounds arbitrary, but it's necessary in order
  // to make shift keys work in a natural way.
  //
  //   The trick is to XOR the current key state with the last key state - the
  // result is a mask with 1 bits where ever a key has changed state.  Then
  // apply the XOR mask to the new state and the result will have a 1 bit only
  // where a key is down now and wasn't down before.  Neat, no?
  //
  //  Lastly, notice that key_press is registered so that it will not actually
  // be asserted until the _next_ clock cycle.  That's the same cycle in which
  // the key output will be updated which is important because we don't want
  // the key_pressed strobe to occur before the data is there!
  wire new_key = key_valid & |(key3 & (keys ^ key3));
  always @(posedge clock)
    key_press <= new_key;
endmodule // ume2_keypad


module ume2_switch_register
  //++
  //   This module implements the DP-8/HM6120 switch register and, as a
  // consequence, manages the two seven segment LED displays.  The UME2
  // displays are used in two distinct modes.  In normal, register display,
  // mode the upper display shows a five digit address in octal (e.g. " 01234")
  // and the lower display shows a single digit register number on the left and
  // a four digit octal value on the right (e.g. "1 4321").  In this mode the
  // register number shows which register's data is being displayed (in other
  // words, it shows us the position of the rotary switch).
  //
  //   The other display mode is used when data is being entered into the switch
  // register.  You enter this mode by pressing any of the number keys, 0-7, and
  // the upper (address) display will blank and the lower (data) display will
  // show the current switch register contents in the format " 0000 ".  Switch
  // register display mode times out after five seconds with no key press, or
  // as soon as any non-numeric key is pressed (e.g. EXAM, LA, LXA, etc).
  //--
#(
  parameter CLOCK_FREQUENCY = 50_000_000,
  parameter DISPLAY_TIMEOUT = 3
) (
  input 	      clock,	// free running 50Mhz system clock
  // FP6120 connections ...
  input [`WORD]       data_leds,// data display LEDs
  input [`WORD]       addr_leds,// address display LEDs
  input [`EMA] 	      ema_leds,	// EMA display LEDs
  input [`ROTSW_BUS]  rotsw,	// current rotary switch setting
  output reg [`WORD]  swreg,	// switch register
  // UME2 keypad and LED connectsions ...
  input  [15:0]	      key,	// current key(s) pressed
  input               key_press,// TRUE for one tick when a key is pressed
  output [6:0] 	      adisp,	// address (upper) 7 segment LEDs segment drive
  output [6:0] 	      ddisp,	// data    (lower) "   "   "   "   "   "    "
  input  [5:0] 	      scan_n	// column strobes for the display
);
`include "clog2.v"

  // Locals ...
  localparam TIMEOUT = CLOCK_FREQUENCY * DISPLAY_TIMEOUT;
  localparam NBITS = clog2(TIMEOUT);
  reg [NBITS-1:0] counter;
  
  function [3:0] RotSwToReg (input [`ROTSW_BUS] rotsw);
  //++
  // Encode the rotary switch position into a register number for display ...
  //--
  begin
    case (rotsw)
      5'b00001: RotSwToReg = 7;		// POST
      5'b00010: RotSwToReg = 1;		// FLAGS
      5'b00100: RotSwToReg = 2;		// AC
      5'b01000: RotSwToReg = 3;		// MQ
      5'b10000: RotSwToReg = 0;		// MD
      default:  RotSwToReg = 4'hF;
    endcase // case (rotsw)
  end
  endfunction // RotSwToReg

  function [2:0] KeyToOctal (input [15:0] key);
  //++
  // Encode a keypad key to it's octal value ...
  //--
  begin
    case (key)
      `KEY_0:  KeyToOctal = 3'o0;
      `KEY_1:  KeyToOctal = 3'o1;
      `KEY_2:  KeyToOctal = 3'o2;
      `KEY_3:  KeyToOctal = 3'o3;
      `KEY_4:  KeyToOctal = 3'o4;
      `KEY_5:  KeyToOctal = 3'o5;
      `KEY_6:  KeyToOctal = 3'o6;
      `KEY_7:  KeyToOctal = 3'o7;
      default: KeyToOctal = 3'o0;
    endcase // case (key)
  end
  endfunction // KeyToOctal

  // TRUE if the current key is any of the number keys ...
  wire is_digit = (key == `KEY_0) | (key == `KEY_1) | (key == `KEY_2)
		| (key == `KEY_3) | (key == `KEY_4) | (key == `KEY_5)
  		| (key == `KEY_6) | (key == `KEY_7);

  // Initialize all registers ...
  initial begin
    swreg = 12'o0000;  counter = 0;
  end
  
  //   This generates the actual switch register.  It's fairly trivial - any
  // time a number key is pressed, the SR shifts left 3 bits and a new digit
  // is added on the right.  The current SR contents are just the last four
  // octal digits entered.  That's all there is to it...
  // Switch register ...
  always @(posedge clock)
    if (key_press & is_digit)
      swreg <= {swreg[3:11], KeyToOctal(key)};

  //   And this generates the display mode timer.  It runs for five full seconds
  // (which is a huge, long time by our standards!) and is started by pressing
  // any numeric key.  It's cleared early by pressing any non-numeric key.
  // The display is in the alternate, switch register display, mode any time
  // the timer is non-zero...
  always @(posedge clock)
    if (key_press)
      counter <= is_digit ? TIMEOUT-1 : 0;
    else if (counter != 0)
      counter <= counter-1;
  wire sw_disp_mode = counter != 0;
  
  //   And lastly generate the drivers for the seven segment displays.  It's
  // pretty easy except for all the multiplexing that goes on to select the
  // appropriate display for the mode ...
  ume2_display #(.ALLOW_HEX(0)) display (
    .adisp(adisp), .ddisp(ddisp), .scan_n(scan_n),
    .addr(sw_disp_mode
            ?  24'hFFFFFF
            : {  4'hF                  , {1'b0, ema_leds},
	        {1'b0, addr_leds[0:2 ]}, {1'b0, addr_leds[3:5 ]},
	        {1'b0, addr_leds[6:8 ]}, {1'b0, addr_leds[9:11]}  }
          ),
    .data(sw_disp_mode
	    ? {  4'hF                  , {1'b0, swreg[0:2 ]},
	        {1'b0, swreg[3:5 ]}    , {1'b0, swreg[6:8 ]},
	        {1'b0, swreg[9:11]}    ,  4'hF                    }
	    : {  RotSwToReg(rotsw)     ,  4'hF, 
	        {1'b0, data_leds[0:2 ]}, {1'b0, data_leds[3:5 ]}, 
	        {1'b0, data_leds[6:8 ]}, {1'b0, data_leds[9:11]}  }
	 )
  );
endmodule // ume2_switch_register


module ume2_ui 
  //++
  //--
#(
  parameter CLOCK_FREQUENCY = 50_000_000
) (
  input 	      clock,	// free running 50Mhz system clock
  // FP6120 connections ...
  input [`WORD]       data_leds,// data display LEDs
  input [`WORD]       addr_leds,// address display LEDs
  input [`EMA] 	      ema_leds,	// EMA display LEDs
  input 	      run_led,	// RUN LED
  input 	      power_led,// POWER LED
  output [`FNSW_BUS]  fnsw,	// function switches (9 of them)
  output reg [`ROTSW_BUS] rotsw,// rotary switch setting
  output [`WORD]  swreg,	// switch register
  // UME2 keypad and LED connectsions ...
  output [6:0] 	      adisp,	// address (upper) 7 segment LEDs segment drive
  output [6:0] 	      ddisp,	// data    (lower) "   "   "   "   "   "    "
  output [5:0] 	      scan_n,	// 7 segment LEDs and keypad column drive
  input  [3:0] 	      keyrow_n,	// keypad row inputs
  output [1:0] 	      led_n,	// two discrete LEDs 
  input  [1:0] 	      sw_n	// two discrete switches
);

  // Create the scan clock and column drivers ....
  wire key_tick;
  ume2_scanner #(.CLOCK_FREQUENCY(CLOCK_FREQUENCY)) scanner
    (.clock(clock), .scan_n(scan_n), .key_tick(key_tick));

  // Keypad scanner ...
  wire [15:0] key;  wire key_press;
  ume2_keypad keypad (
    .clock(clock), .scan_n(scan_n), .key_tick(key_tick),
    .keyrow_n(keyrow_n), .keys(key), .key_press(key_press)
  );

  ume2_switch_register #(.CLOCK_FREQUENCY(CLOCK_FREQUENCY)) sr (
    .clock(clock), .data_leds(data_leds), .addr_leds(addr_leds),
    .ema_leds(ema_leds), .rotsw(rotsw), .swreg(swreg), .key(key),
    .key_press(key_press), .adisp(adisp), .ddisp(ddisp), .scan_n(scan_n)
  );

  // Rotary switch ...
  initial rotsw = 5'b10000;
  always @(posedge clock)
         if (key_press & (key == `KEY_MD))
      rotsw <= 5'b10000;
    else if (key_press & (key == `KEY_FLAGS))
      rotsw <= 5'b00010;
    else if (key_press & (key == `KEY_AC))
      rotsw <= 5'b00100;
    else if (key_press & (key == `KEY_MQ))
      rotsw <= 5'b01000;
    else if (key_press & (key == `KEY_POST))
      rotsw <= 5'b00001;
    
  assign fnsw[`FNSW_LA]    = key == `KEY_LA;
  assign fnsw[`FNSW_LXA]   = key == `KEY_LXA;
  assign fnsw[`FNSW_EXAM]  = key == `KEY_EXAM;
  assign fnsw[`FNSW_DEP]   = key == `KEY_DEP;
  assign fnsw[`FNSW_CLEAR] = key == `KEY_CLEAR;
  assign fnsw[`FNSW_CONT]  = key == `KEY_CONT;
  assign fnsw[`FNSW_BOOT]  = key == `KEY_BOOT;

  wire sw_halt, sw_lock;
  debouncer #(.ACTIVE_STATE(0))
    halt_debounce (.clock(clock), .switch(sw_n[0]), .state(sw_halt) );
  debouncer #(.ACTIVE_STATE(0))
    lock_debounce (.clock(clock), .switch(sw_n[1]), .state(sw_lock) );
  assign fnsw[`FNSW_LOCK] = sw_lock;
  assign fnsw[`FNSW_HALT] = sw_halt;

  // Two of the UME2 LEDs are used for the POWER and RUN LEDs ...  
  assign led_n[0] = ~power_led;
  assign led_n[1] = ~run_led;
endmodule // ume2_ui


module sbc6120_ume2 (
  // S3 board I/Os from s2.ucf ....
  input        clock_50mhz_in,	// 50MHz master clock
//output       slu0_txd,	// RS232/female DB9 TXD
//input        slu0_rxd,	// RS232/female DB9 RXD
  // SRAM connections ...
  output [18:0]ram_ma,		// SRAM address bits
  inout  [11:0]ram_md,		// SRAM data bits
  output       ram_oe_n,	// SRAM output enable
  output       ram_we_high_n,	// SRAM write enable (high byte)
  output       ram_we_low_n,	// SRAM write enable (low byte)
  // PS/2 keyboard connections ...
  inout	       ps2_clock_n,	// PS/2 keyboard clock
  inout	       ps2_data_n,	// PS/2 keyboard data
  // VGA connections ...
  output       vga_red,		// VGA red video
  output       vga_green,	// VGA green video
  output       vga_blue,	// VGA blue video
  output       vga_hsync,	// VGA horizontal sync
  output       vga_vsync,	// VGA vertical sync
  // CompactFlash card interface (in common memory model mode) ...
  output [2:0] cf_a,		// register select bits
  inout  [7:0] cf_d,		// 8 bit data bus
  output       cf_oe_n,		// output enable (read strobe)
  output       cf_we_n,		// write strobe
  output       cf_cs_n,		// card select
  output       cf_reset,	// reset the card
  input        cf_ready_n,	// card ready
  input        cf_cd_n,		// card inserted
  // MMC/SD card SPI interface ...
  output       mmc_sclk,	// SPI clock
  output       mmc_mosi,	// master (that's us!) our, slave in
  input        mmc_miso,	// master in, slave out
  output       mmc_cs_n,	// slave select
  input        mmc_cd_n,	// card detected
  input        mmc_wp_n,	// card is write protectedz
  // DS1302 interface ...
  output       rtc_sclk,	// serial clock
  output       rtc_ce,		// chip enable and byte sync
  inout	       rtc_sio,		// bidirectional serial data
  // UME2 keypad and LED connectsions ...
  output [6:0] adisp,		// address (upper) 7 segment LEDs segment drive
  output [6:0] ddisp,		// data    (lower) "   "   "   "   "   "    "
  output [5:0] scan_n,		// 7 segment LEDs and keypad column drive
  input  [3:0] keyrow_n,	// keypad row inputs
  output [1:0] led_n,		// two LEDs (UME2 has four, but we only use two)
  input  [1:0] sw_n,		// two switches (again, out of four)
  output       speaker,		// push pull drive for the piezo beeper
  output       speaker_n	// ...
);
  // Parameters ...
  parameter CLOCK_FREQUENCY      = 50_000_000;
  parameter CPU_CLOCK_DIVIDE     = 4;
  parameter CONSOLE_BAUD_RATE    = 19200;
  parameter PIXEL_CLOCK_MULTIPLY = 17;
  parameter PIXEL_CLOCK_DIVIDE   = 30;
  localparam CPU_CLOCK_FREQUENCY = CLOCK_FREQUENCY / CPU_CLOCK_DIVIDE;
  localparam PIXEL_FREQUENCY     = (CLOCK_FREQUENCY * PIXEL_CLOCK_MULTIPLY) / PIXEL_CLOCK_DIVIDE;

  // Locals ... 
  wire clock_50mhz_buf, vgaclk, cpuclk;
  wire sbc6120_txd, sbc6120_rxd, vt52_txd, vt52_rxd, bell;
  wire [2:0] post_leds;
`ifdef FP6120
  wire run_led, power_led;
  wire [`WORD] data_leds, addr_leds, swreg;  wire [`EMA] ema_leds;
  wire [`FNSW_BUS] fnsw;  wire [`ROTSW_BUS] rotsw;
`endif
`ifdef XRAM
  wire ram_we_n;
`endif
 
  // Clocks ...
  IBUFG clock_50mhz_ibufg (.I(clock_50mhz_in), .O(clock_50mhz_buf));
  ume2_clkgen #(
    .CPU_CLOCK_DIVIDE(CPU_CLOCK_DIVIDE),
    .PIXEL_CLOCK_MULTIPLY(PIXEL_CLOCK_MULTIPLY),
    .PIXEL_CLOCK_DIVIDE(PIXEL_CLOCK_DIVIDE)
  ) ume2_clkgen (
    .clock_50mhz(clock_50mhz_buf), .cpuclk(cpuclk), .vgaclk(vgaclk)
  );
    
  // Here's the important part... 
  sbc6120 #(
    .CPU_CLOCK(CPU_CLOCK_FREQUENCY), .CONSOLE_BAUD(CONSOLE_BAUD_RATE)
  ) sbc6120 (
    .cpuclk(cpuclk), .post_code(post_leds),
`ifdef XRAM
    .xram_ma(ram_ma[15:0]), .xram_md(ram_md[11:0]),
    .xram_oe_n(ram_oe_n), .xram_we_n(ram_we_n),
`endif
`ifdef CFCARD
    .cf_a(cf_a), .cf_d(cf_d), .cf_oe_n(cf_oe_n), .cf_we_n(cf_we_n),
    .cf_cd_n(cf_cd_n), .cf_cs_n(cf_cs_n), .cf_reset(cf_reset),
    .cf_ready_n(cf_ready_n),
`endif
`ifdef SDCARD
    .mmc_sclk(mmc_sclk), .mmc_mosi(mmc_mosi), .mmc_miso(mmc_miso),
    .mmc_cs_n(mmc_cs_n), .mmc_cd_n(mmc_cd_n), .mmc_wp_n(mmc_wp_n),
`endif
`ifdef RTC
    .rtc_sclk(rtc_sclk), .rtc_ce(rtc_ce), .rtc_sio(rtc_sio),
`endif
`ifdef FP6120
    .data_leds(data_leds), .addr_leds(addr_leds), .ema_leds(ema_leds),
    .run_led(run_led), .power_led(power_led),
    .swreg(swreg), .fnsw(fnsw), .rotsw(rotsw),
`endif
    .console_rxd(sbc6120_rxd), .console_txd(sbc6120_txd)
  );

  // XRAM interface
`ifdef XRAM
  assign ram_we_high_n = ram_we_n;  assign ram_we_low_n = ram_we_n;
  assign ram_ma[18:16] = 3'b0;  //assign ram_md[15:12] = 4'bz;
`else  
  assign ram_we_high_n = 1'b1;  assign ram_we_low_n = 1'b1;
  assign ram_oe_n = 1'b1;
  assign ram_ma = 19'b0;  assign ram_md = 15'b0;
`endif // !`ifdef XRAM

  //   The CPU and VT52 have separate clock domains (cpuclk vs vgaclk, of
  // course) and there are exactly two signals that cross between them - TXD
  // and RXD.  This creates synchronizers for those two signals.  That's
  // probably not really necessary, but it seems like a good idea...
  synchronize_level cpu2vga (.clock(vgaclk), .in(sbc6120_txd), .out(vt52_rxd));
  synchronize_level vga2cpu (.clock(cpuclk), .in(vt52_txd), .out(sbc6120_rxd));

  // VT52 console terminal...
  vt52 #(
    .CLOCK_FREQUENCY(PIXEL_FREQUENCY), .BAUD_RATE(CONSOLE_BAUD_RATE),
    .FOREGROUND(`RGB_YELLOW), .BACKGROUND(`RGB_BLACK),
    .CURS_BLINK(1'b1), .CURS_UNDERLINE(1'b0), .AUTO_NEWLINE(1'b1),
    .MARGIN_BELL(1'b1), .SWAP_CAPS_CTRL(1'b1), .INIT_KEYPAD_MODE(1'b0),
    .RESET_KEYBOARD(1'b1)
  ) vt52 (
    .clock(vgaclk), .rxd(vt52_rxd), .txd(vt52_txd),
    .ps2_clock(ps2_clock_n), .ps2_data(ps2_data_n),
    .hsync(vga_hsync), .vsync(vga_vsync), .bell(bell),
    .video({vga_red, vga_green, vga_blue})
  );
  ume2_beeper beeper (
    .clock(vgaclk), .enable(bell), .speaker(speaker), .speaker_n(speaker_n)
  );

 // User interface (aka the "front panel") ...
`ifdef FP6120
  ume2_ui #(.CLOCK_FREQUENCY(CPU_CLOCK_FREQUENCY)) ui (
    .clock(cpuclk), .swreg(swreg),
    .data_leds(data_leds), .addr_leds(addr_leds), .ema_leds(ema_leds),
    .run_led(run_led), .power_led(power_led), .fnsw(fnsw), .rotsw(rotsw),
    .adisp(adisp), .ddisp(ddisp), .scan_n(scan_n),
    .keyrow_n(keyrow_n), .led_n(led_n), .sw_n(sw_n)
  );
`endif

  // Disable CF card when no interface is generated ...
`ifndef CFCARD
  assign cf_a = 3'b0;  assign cf_d = 8'b0;  assign cf_reset = 1'b0;
  assign cf_oe_n = 1'b1;  assign cf_we_n = 1'b1;  assign cf_cs_n = 1'b1;
`endif
  // Disable MMC/SD card when no interface is generated ...
`ifndef SDCARD
  assign mmc_sclk = 1'b0;  assign mmc_mosi = 1'b0;  assign mmc_cs_n = 1'b1;
`endif
  // Disable DS1302 when no interface is generated ...
`ifndef RTC
  assign rtc_sclk = 1'b0;  assign rtc_ce = 1'b0;  assign rtc_sio = 1'b0;
`endif
  // Disable UME2 LEDs when no FP6120 is generated ...
`ifndef FP6120
  assign adisp = 7'h00;  assign ddisp = 7'h00;  assign scan_n = 6'h3F;
  assign led_n = {1'b1, 1'b1};
`endif

endmodule // sbc6120_ume2
