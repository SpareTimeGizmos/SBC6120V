//++
//sbc6120_s3.v
//
//   SBC6120V TEST BENCH FOR DIGILENT S3 STARTER BOARD
//   Copyright (C) 2011 by Spare Time Gizmos.  All rights reserved.
//
// DESIGN NAME:	SBC6120V
// DESCRIPTION:
//   This module runs the SBC6120V on the Digilent S3 evaluation board.  The
// actual FPGA on the board I used is the Spartan 3 XC3S400-5ft256 - there
// are other versions of the board with XC3S200 and XC3S1000 parts that would
// probably work equally well.
//
// The S3 board has no CompactFlash interface and no mass storage.  Sorry.
//
// Be sure to use the S3.UCF constrants file when building this design!
//
// Currently this design uses the 8 discrete LEDs as follows-
//
//	LED 7 - RESET
//	LED 6 - console activity (TXD or RXD)
//	LED 5 - visible "bell"
//	LED 4 - unused
//	LED 3 - always on (like the POWER led on the SBC6120)
//	LED 2 - POST code (MSB)
//	LED 1 - POST code
//	LED 0 - POST code (LSB)
//
// Push button 3 is a reset, as is common with many S3 designs.
//
// The remaining push buttons, the eight slide switches, and the seven
// segment display are currently unused.
//
// REVISION HISTORY:
// 22-Jan-11 RLA  new file.
//--
//000000011111111112222222222333333333344444444445555555555666666666677777777778
//345678901234567890123456789012345678901234567890123456789012345678901234567890
`include "sbc6120_h.v"


module s3_clkgen
  //++
  //   This module uses one of the nifty Xilinx digital clock managers to
  // generate both a CPU clock and a VGA pixel clock.  The system clock is
  // nominally 50Mhz and a 25MHz CPU clock is generated by using the DLL part
  // of the DCM to divide by two.  At the same time we use the frequency
  // synthesizer part of the same DCM to generate a 28.322MHz VGA dot clock
  // by multiplying the ratio 17/30.  That's all there is to it!
  //--
( 
  input  clock_50mhz, 	// 50Mhz system clock
  output cpuclk, 	// 25Mhz cpu clock
  output vgaclk,	// 28.322Mhz VGA dot clock
  output locked		// TRUE when the DCM is locked
);
  parameter CPU_CLOCK_DIVIDE     =  2;
  parameter PIXEL_CLOCK_MULTIPLY = 17;
  parameter PIXEL_CLOCK_DIVIDE   = 30;

  // Locals ...
  wire clkdv_unbuf;	// unbuffered DCM CLKDV (cpuclk)
  wire clkfx_unbuf;	// unbuffered DCM CLKFX (vgaclk)
  wire clk0_unbuf;	// unbuffered DCM CLK0 output
  wire clkfb_buf;	// buffered CLK0 for DCM feedback

  // Here's the magic part!
  DCM #(
    .CLKDV_DIVIDE(CPU_CLOCK_DIVIDE),
    .CLKFX_DIVIDE(PIXEL_CLOCK_DIVIDE), .CLKFX_MULTIPLY(PIXEL_CLOCK_MULTIPLY),
    .CLK_FEEDBACK("1X"), .FACTORY_JF(16'h8080)
   ) clkdcm (
    .CLKIN(clock_50mhz), .CLK0(clk0_unbuf), .CLKFB(clkfb_buf), 
    .CLKDV(clkdv_unbuf), .CLKFX(clkfx_unbuf), .LOCKED(locked),
    .DSSEN(0), .PSCLK(0), .PSEN(0), .PSINCDEC(0), .RST(0)
  );
  
  //   Buffer all the clocks we generate with global buffers, and that includes
  // sticking a BUFG in the feedback path for the DCM.  That's so the DCM will
  // automatically compensate for the 1ns or so delay added by the BUFG.  This
  // application is not very critical and that's overkill, but it's the "right" 
  // way to do it...
  BUFG cpuclk_bufg    (.I(clkdv_unbuf), .O(cpuclk));
  BUFG vgaclk_bufg    (.I(clkfx_unbuf), .O(vgaclk));
  BUFG clkdcm_fb_bufg (.I(clk0_unbuf),  .O(clkfb_buf));
endmodule // s3_clkgen


module s3_reset
  //++
  //   This module implements the logic for resetting the SBC6120.  It's
  // primary purpose is to hold the system in the reset state until all DCMs
  // have locked and stayed locked for at least 50ms.  Yes, 50ms is a huge
  // long time but we don't really care.
  //
  //   It's secondary purpose is to hold reset asserted for at least 50ms
  // after the reset push button is pressed.  In this application the long
  // timeout is handy because it means we don't need any other debouncing
  // for the button...
  //--
(
  input  sysclk,	// free running 50Mhz system clock
  input  locked,	// all DCMs have locked
  input  button,	// external reset push button
  output reset		// system reset
);
  parameter LOG2_DELAY = 22;
  reg [LOG2_DELAY-1:0] count;

  always @(posedge sysclk)
    if (button | !locked)
      count <= 2**LOG2_DELAY-1;
    else if (count != 0)
      count <= count - 1;
      
  assign reset = count != 0;
endmodule // s3_reset


module s3_bell (
  //   This module is supposed to ring the bell, however the S3 board doesnt'
  // have one.  We'll just fake it by blinking an LED instead...
  //--
  input  sysclk,	// free running 50Mhz system clock
  input  reset,		// global asynchronous reset
  input  bell,		// asserted for one tick to trigger the bell
  output led		// drive an LED with this
);
  parameter LOG2_DELAY = 23; // about 0.16s at 50Mhz
  reg [LOG2_DELAY-1:0] count;
  
  always @(posedge sysclk or posedge reset)
    if (reset)
      count <= 0;
    else if (bell)
      count <= 2**LOG2_DELAY-1;
    else if (count != 0)
      count <= count-1;
 
  assign led = count != 0;
endmodule // s3_bell


module sbc6120_s3 (
  // S3 board I/Os from s2.ucf ....
  input        clock_50mhz_in,	// 50MHz master clock
  input        reset_button,	// reset push button
  output [7:0] leds,		// discrete LEDs (not the 7 segment display!)
//output       txd,		// RS232/female DB9 TXD
//input        rxd,		// RS232/female DB9 RXD
  output [17:0]ram_addr,	// SRAM address bits
  output       ram_oe_n,	// SRAM output enable
  output       ram_we_n,	// SRAM write enable
  inout  [11:0]ram_a_data,	// SRAM "a" data
  output       ram_a_ce_n,	// SRAM "a" chip enable
  output       ram_a_lb_n,	// SRAM "a" lower byte enable
  output       ram_a_ub_n,	// SRAM "a" upper byte enable
//inout  [15:0]ram_b_data,	// SRAM "b" data
  output       ram_b_ce_n,	// SRAM "b" chip enable
  output       ram_b_lb_n,	// SRAM "b" lower byte enable
  output       ram_b_ub_n,	// SRAM "b" upper byte enable
  inout	       ps2_clock,	// PS/2 keyboard clock
  inout	       ps2_data,	// PS/2 keyboard data
  output       vga_red,		// VGA red video
  output       vga_green,	// VGA green video
  output       vga_blue,	// VGA blue video
  output       vga_hsync,	// VGA horizontal sync
  output       vga_vsync	// VGA vertical sync
//input	[2:0] btn		// temporary!!
);
  parameter CLOCK_FREQUENCY      = 50_000_000;
  parameter CPU_CLOCK_DIVIDE     = 2;
  parameter CONSOLE_BAUD_RATE    = 19200;
  parameter PIXEL_CLOCK_MULTIPLY = 17;
  parameter PIXEL_CLOCK_DIVIDE   = 30;
  localparam CPU_CLOCK_FREQUENCY = CLOCK_FREQUENCY / CPU_CLOCK_DIVIDE;
  localparam PIXEL_FREQUENCY     = (CLOCK_FREQUENCY * PIXEL_CLOCK_MULTIPLY) / PIXEL_CLOCK_DIVIDE;
  
  // Clocks ...
  wire clkdcm_locked, clock_50mhz_buf, vgaclk, cpuclk;
  IBUFG clock_50mhz_ibufg (.I(clock_50mhz_in), .O(clock_50mhz_buf));
  s3_clkgen #(
    .CPU_CLOCK_DIVIDE(CPU_CLOCK_DIVIDE),
    .PIXEL_CLOCK_MULTIPLY(PIXEL_CLOCK_MULTIPLY),
    .PIXEL_CLOCK_DIVIDE(PIXEL_CLOCK_DIVIDE)
  ) s3_clkgen (
    .clock_50mhz(clock_50mhz_buf), .locked(clkdcm_locked),
    .cpuclk(cpuclk), .vgaclk(vgaclk)
  );
    
  // Reset logic ...  
  wire reset;
  s3_reset #(24) s3_reset (
    .sysclk(clock_50mhz_buf), .button(reset_button),
    .locked(clkdcm_locked), .reset(reset)
  );

  // Here's the important part... 
  wire console_txd, console_rxd;
  sbc6120 #(
    .CPU_CLOCK(CPU_CLOCK_FREQUENCY),
    .CONSOLE_BAUD(CONSOLE_BAUD_RATE)
  ) sbc6120 (
    .cpuclk(cpuclk), .reset(reset), .leds(leds[2:0]),
    .xram_ma(ram_addr[15:0]), .xram_md(ram_a_data[11:0]),
    .xram_oe_n(ram_oe_n), .xram_we_n(ram_we_n),
    .ide_da(), .ide_dd(), .ide_dior_n(), .ide_diow_n(),
    .ide_cs1fx_n(), .ide_cs3fx_n(), .ide_dreset_n(), .ide_dasp_n(0),
    .console_rxd(console_rxd), .console_txd(console_txd)
  );
  
  // RAM "a" is always selected and RAM "b" is disabled ...
  assign ram_a_ce_n = 0;  assign ram_a_lb_n = 0;  assign ram_a_ub_n = 0;
  assign ram_b_ce_n = 1;  assign ram_b_lb_n = 1;  assign ram_b_ub_n = 1;
  assign ram_addr[17:16] = 2'b0;  //assign ram_a_data[15:12] = 4'bz;

  wire bell;
  vt52 #(
    .CLOCK_FREQUENCY(PIXEL_FREQUENCY),
    .BAUD_RATE(CONSOLE_BAUD_RATE),
    .FOREGROUND(`RGB_YELLOW),
    .BACKGROUND(`RGB_BLACK),
    .CURS_BLINK(1),
    .CURS_UNDERLINE(0),
    .AUTO_NEWLINE(1),
    .MARGIN_BELL(1),
    .SWAP_CAPS_CTRL(1),
    .INIT_KEYPAD_MODE(0),
    .RESET_KEYBOARD(1)
  ) vt52 (
    .clock(vgaclk), .reset(reset),
    .rxd(console_txd), .txd(console_rxd),
    .ps2_clock(ps2_clock), .ps2_data(ps2_data),
    .hsync(vga_hsync), .vsync(vga_vsync), .video({vga_blue, vga_green, vga_red}),
    .bell(bell)
  );
  s3_bell s3_bell (
    .sysclk(vgaclk), .reset(reset), .bell(bell), .led(leds[5])
  );

  // Drive the LEDs on the S3 board...
  assign leds[4] = 0;  assign leds[3] = 1;
  assign leds[7] = reset;
  assign leds[6] = (~console_txd) | (~console_rxd);
endmodule

